`ifndef NOTE_TABLE_VH
`define NOTE_TABLE_VH

`define NOTE_RST  6'd0    //     0.00000 Hz

`define NOTE_A2   6'd1    //   110.00000 Hz

`define NOTE_C3   6'd2    //   130.81280 Hz
`define NOTE_D3   6'd3    //   146.83240 Hz
`define NOTE_Ds3  6'd4    //   155.56350 Hz
`define NOTE_E3   6'd5    //   164.81380 Hz
`define NOTE_F3   6'd6    //   174.61410 Hz
`define NOTE_Fs3  6'd7    //   184.99720 Hz
`define NOTE_G3   6'd8    //   195.99770 Hz
`define NOTE_A3   6'd9    //   220.00000 Hz
`define NOTE_As3  6'd10   //   233.08190 Hz
`define NOTE_B3   6'd11   //   246.94170 Hz

`define NOTE_C4   6'd12   //   261.62560 Hz
`define NOTE_Cs4  6'd13   //   277.18260 Hz
`define NOTE_D4   6'd14   //   293.66480 Hz
`define NOTE_Ds4  6'd15   //   311.12700 Hz
`define NOTE_E4   6'd16   //   329.62760 Hz
`define NOTE_F4   6'd17   //   349.22820 Hz
`define NOTE_Fs4  6'd18   //   369.99440 Hz
`define NOTE_Gs4  6'd19   //   415.30470 Hz
`define NOTE_A4   6'd20   //   440.00000 Hz
`define NOTE_As4  6'd21   //   466.16380 Hz
`define NOTE_B4   6'd22   //   493.88330 Hz

`define NOTE_C5   6'd23   //   523.25110 Hz
`define NOTE_Cs5  6'd24   //   554.36530 Hz
`define NOTE_Fs5  6'd25   //   739.98880 Hz
`define NOTE_Gs5  6'd26   //   830.60940 Hz
`define NOTE_A5   6'd27   //   880.00000 Hz
`define NOTE_As5  6'd28   //   932.32750 Hz
`define NOTE_B5   6'd29   //   987.76660 Hz

`define NOTE_C6   6'd30   //  1046.50200 Hz
`define NOTE_Cs6  6'd31   //  1108.73100 Hz
`define NOTE_Fs6  6'd32   //  1479.97800 Hz
`define NOTE_Gs6  6'd33   //  1661.21900 Hz
`define NOTE_A6   6'd34   //  1760.00000 Hz
`define NOTE_As6  6'd35   //  1864.65500 Hz
`define NOTE_B6   6'd36   //  1975.53300 Hz

`define NOTE_Cs7  6'd37   //  2217.46100 Hz

`endif
