`ifndef NOTE_TABLE_VH
`define NOTE_TABLE_VH

`define NOTE_RST  6'd0    //     0.00000 Hz

`define NOTE_A1   6'd1    //   110.00000 Hz

`define NOTE_C2   6'd2    //   130.81280 Hz
`define NOTE_D2   6'd3    //   146.83240 Hz
`define NOTE_E2   6'd4    //   164.81380 Hz
`define NOTE_F2   6'd5    //   174.61410 Hz
`define NOTE_Fs2  6'd6    //   184.99720 Hz
`define NOTE_G2   6'd7    //   195.99770 Hz
`define NOTE_A2   6'd8    //   220.00000 Hz
`define NOTE_B2   6'd9    //   246.94170 Hz

`define NOTE_C3   6'd10   //   261.62560 Hz
`define NOTE_Cs3  6'd11   //   277.18260 Hz
`define NOTE_D3   6'd12   //   293.66480 Hz
`define NOTE_E3   6'd13   //   329.62760 Hz
`define NOTE_F3   6'd14   //   349.22820 Hz
`define NOTE_Fs3  6'd15   //   369.99440 Hz
`define NOTE_Gs3  6'd16   //   415.30470 Hz
`define NOTE_A3   6'd17   //   440.00000 Hz
`define NOTE_As3  6'd18   //   466.16380 Hz
`define NOTE_B3   6'd19   //   493.88330 Hz

`define NOTE_C4   6'd20   //   523.25110 Hz
`define NOTE_Cs4  6'd21   //   554.36530 Hz
`define NOTE_Fs4  6'd22   //   739.98880 Hz
`define NOTE_Gs4  6'd23   //   830.60940 Hz
`define NOTE_A4   6'd24   //   880.00000 Hz
`define NOTE_As4  6'd25   //   932.32750 Hz
`define NOTE_B4   6'd26   //   987.76660 Hz

`define NOTE_C5   6'd27   //  1046.50200 Hz
`define NOTE_Cs5  6'd28   //  1108.73100 Hz
`define NOTE_Fs5  6'd29   //  1479.97800 Hz
`define NOTE_Gs5  6'd30   //  1661.21900 Hz
`define NOTE_A5   6'd31   //  1760.00000 Hz
`define NOTE_As5  6'd32   //  1864.65500 Hz
`define NOTE_B5   6'd33   //  1975.53300 Hz

`define NOTE_Cs6  6'd34   //  2217.46100 Hz

`endif
