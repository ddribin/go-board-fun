`ifndef _NES_CONTROLLER_VH
`define _NES_CONTROLLER_VH

`define NES_BUTTON_A      3'd7
`define NES_BUTTON_B      3'd6
`define NES_BUTTON_SELECT 3'd5
`define NES_BUTTON_START  3'd4
`define NES_BUTTON_UP     3'd3
`define NES_BUTTON_DOWN   3'd2
`define NES_BUTTON_LEFT   3'd1
`define NES_BUTTON_RIGHT  3'd0

`endif
