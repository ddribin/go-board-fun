module pwm_top (
);
  
endmodule
