`ifndef NOTE_TABLE_VH
`define NOTE_TABLE_VH

`define NOTE_RST  6'd0    //     0.00000 Hz

`define NOTE_A2   6'd1    //   110.00000 Hz

`define NOTE_C3   6'd2    //   130.81280 Hz
`define NOTE_D3   6'd3    //   146.83240 Hz
`define NOTE_E3   6'd4    //   164.81380 Hz
`define NOTE_F3   6'd5    //   174.61410 Hz
`define NOTE_G3   6'd6    //   195.99770 Hz
`define NOTE_A3   6'd7    //   220.00000 Hz
`define NOTE_B3   6'd8    //   246.94170 Hz

`define NOTE_C4   6'd9    //   261.62560 Hz
`define NOTE_D4   6'd10   //   293.66480 Hz
`define NOTE_E4   6'd11   //   329.62760 Hz
`define NOTE_F4   6'd12   //   349.22820 Hz
`define NOTE_Fs4  6'd13   //   369.99440 Hz
`define NOTE_A4   6'd14   //   440.00000 Hz

`define NOTE_C5   6'd15   //   523.25110 Hz
`define NOTE_Cs5  6'd16   //   554.36530 Hz
`define NOTE_Fs5  6'd17   //   739.98880 Hz
`define NOTE_Gs5  6'd18   //   830.60940 Hz
`define NOTE_A5   6'd19   //   880.00000 Hz
`define NOTE_As5  6'd20   //   932.32750 Hz
`define NOTE_B5   6'd21   //   987.76660 Hz

`endif
