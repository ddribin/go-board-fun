`default_nettype none
module nes_controller #(
  clk_freq_hz = 0
) (
  input wire      i_clk,
  output wire     o
);

  assign o = 1;
  
endmodule
